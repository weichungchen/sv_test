module test
{
    input a;
    output b;
};

    assign b = a + 1'd1;

endmodule
