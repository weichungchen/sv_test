module test
{
    input a;
    output b;
};
endmodule
