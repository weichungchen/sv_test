module test
{
    input a;
    output b;
};

    assign b =  a;

endmodule
